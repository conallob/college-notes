-- $Id: splitter.vhd,v 1.3 2004/04/14 21:52:35 conall Exp $


