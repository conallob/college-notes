library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity 2to1mux is
    Port ( );
end 2to1mux;

architecture Behavioral of 2to1mux is

begin


end Behavioral;
